-------------------------------------------------------------------------------------
-- Transceiver Hardware Component Container, version 2 (for Mk8 Apex/XCVR)
-------------------------------------------------------------------------------------
-- Author:      Maxwell Phillips
-- Copyright:   Ohio Northern University, 2023.
-- License:     GPL v3
-- Description: Container for hardware to be wrapped by apex component.
-------------------------------------------------------------------------------------
--
-- This file is the hardware component container wrapped by the top level apex
-- component. You should modify this file to wrap your hardware in order to utilize
-- it with the serial transceiver. See the apex component and transceiver files
-- for more details on their functionality.
--
-------------------------------------------------------------------------------------
-- Generics
-------------------------------------------------------------------------------------
--
-- [G_byte_bits]: Should be 8. Mapped from top-level component.
--
-- [G_total_bits]: The capacity, in bits, of the transceiver.
--                 Mapped directly from the top-level component.
--                 Should be used to help structure hardware components.
--
-- [G_clk_freq]: Should match the clock frequency of the FPGA board.
--               Again, mapped by top-level component.
--
-------------------------------------------------------------------------------------
-- Ports
-------------------------------------------------------------------------------------
--
-- [clk_100mhz]: Input clock signal; should match [G_clk_freq] generic.
--
-- [clk_hw]: Clock signal to time contained hardware. Generated by MMCM on top-level.
--
-- [reset]: Asynchronous reset signal. The module should be initially
--          reset automatically by the transceiver, and will remain reset
--          until all bytes are received and the processing stage begins.
--          To preserve state, the hardware is NOT reset after the processing
--          stage and during the transmission stage. This allows displaying
--          output on the LEDs from the hardware container more easily.
--
-- [load]: Signal which is received for one clock cycle (of [G_clk_freq]) at the
--         beginning of the processing stage, to allow for any hardware setup.
--
-- [start]: Signal which is asserted for as long as the processing stage is active.
--          Will remain high until [done] is asserted.
--
-- [btn_X]: These four signals are mapped to their corresponding buttons
--          on the FPGA development board. By default, left and right are
--          used by the transceiver to display the delay counter on the LEDs.
--          In order to utilize the LEDs for your hardware, you must assert
--          [override_leds] when a button is pressed and set [leds] as desired.
--
-- [switches]: The 16 dip switches on the FPGA development board.
--
-- [input]: Parallel input of size [G_total_bits] from the transceiver.
--
-- [output]: Parallel output of size [G_total_bits] back to the transceiver.
--
-- [done]: Done signal for the transceiver to terminate the processing stage
--         and begin to transmit the result (from [output]) back over UART.
--
-- [override_leds]: Signal to use [leds] from the hardware instead of transceiver.
--
-- [leds]: Output LEDs. Controlled by the top-level component based on [override_leds].
--
-------------------------------------------------------------------------------------

library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.numeric_std.all;
  use IEEE.std_logic_unsigned.all;
  use IEEE.math_real.all;

entity hw_container is
  generic (
    G_byte_bits  : integer;
    G_total_bits : integer;
    G_clk_freq   : integer
  );
  port (
    clk_100mhz    : in    std_logic; -- board clk
    clk_hw        : in    std_logic; -- clock to be passed to hardware
    reset         : in    std_logic; -- async reset which is high when xcvr is not in processing stage
    load          : in    std_logic; -- pseudo-async pulse received from xcvr at the start of processing stage
    start         : in    std_logic; -- consistent signal received from xcvr as long as processing stage is active
    btn_up        : in    std_logic;
    btn_left      : in    std_logic; -- left is by default used for displaying left half of delay counter from xcvr
    btn_right     : in    std_logic; -- right is by default used for displaying right half of delay counter from xcvr
    btn_down      : in    std_logic;
    switches      : in    std_logic_vector(15 downto 0);
    input         : in    std_logic_vector(G_total_bits - 1 downto 0);
    output        : out   std_logic_vector(G_total_bits - 1 downto 0);
    done          : out   std_logic; -- tells xcvr to finish processing stage and transmit back result ([output])
    override_leds : out   std_logic; -- tells xcvr to use [leds] instead of displaying bytes received or delay
    leds          : out   std_logic_vector(15 downto 0)
  );
end hw_container;

architecture behavioral of hw_container is

  -- divider
  constant G_n : integer := G_total_bits / 2;

  -- don't override generics since this algorithm is not fully generalizable
  component division_algorithm_1024 is
    port (
      clk       : in    std_logic;
      reset     : in    std_logic;
      load      : in    std_logic;
      start     : in    std_logic;
      s_dd      : in    std_logic;
      dividend  : in    std_logic_vector(G_n - 1 downto 0);
      s_dr      : in    std_logic;
      divisor   : in    std_logic_vector(G_n - 1 downto 0);
      done      : out   std_logic;
      s_q       : out   std_logic;
      quotient  : out   std_logic_vector(G_n - 1 downto 0);
      s_r       : out   std_logic;
      remainder : out   std_logic_vector(G_n - 1 downto 0)
    );
  end component;

  -- divider data signals
  signal s_dr   : std_logic;
  signal s_dd   : std_logic;
  signal s_q    : std_logic;
  signal s_r    : std_logic;
  signal mag_dr : std_logic_vector(G_n - 1 downto 0);
  signal mag_dd : std_logic_vector(G_n - 1 downto 0);
  signal mag_q  : std_logic_vector(G_n - 1 downto 0);
  signal mag_r  : std_logic_vector(G_n - 1 downto 0);

  -- divider logistics signals
  signal dr_hw_reset : std_logic;
  signal dr_hw_done  : std_logic;

begin

  s_dd   <= switches(15);
  mag_dd <= input(input'left downto G_n);
  s_dr   <= switches(14);
  mag_dr <= input(G_n - 1 downto 0);

  dr_hw_reset <= reset;
  done        <= dr_hw_done;
  output      <= mag_q & mag_r;

  process (clk_100mhz, reset) begin
    if (reset = '1') then
      override_leds <= '0'; -- IMPORTANT!
      leds          <= (others => '0');
    elsif (clk_100mhz'event and clk_100mhz = '1') then
      -- LED multiplexing
      if (btn_down = '1') then
        override_leds     <= '1';
        leds(15)          <= s_dd;
        leds(14)          <= s_dr;
        leds(13 downto 2) <= (others => '0');
        leds(1)           <= s_q;
        leds(0)           <= s_r;
      else
        override_leds <= '0';
      end if;
    end if;
  end process;

  divider : division_algorithm_1024
    port map (
      clk       => clk_hw,
      reset     => dr_hw_reset,
      load      => load,
      start     => start,
      s_dd      => s_dd,
      dividend  => mag_dd,
      s_dr      => s_dr,
      divisor   => mag_dr,
      done      => dr_hw_done,
      s_q       => s_q,
      quotient  => mag_q,
      s_r       => s_r,
      remainder => mag_r
    );

end architecture behavioral;
